.title TestCircuit
Ra in p1 5
Rb p1 0 5
Vin in 0 DC 9
.op
.print op v(p1)

