.title TestCircuit
Ra vin p1 5
Rb p1 0 5
Vin vin 0 DC 0 EXTERNAL
.op
.print op v(p1)
